.SUBCKT MCP606 1 2 3 4 5
*              | | | | |
*              | | | | Output
*              | | | Negative Supply
*              | | Positive Supply
*              | Inverting Input
*              Non-inverting Input
*
********************************************************************************
* Software License Agreement                                                   *
*                                                                              *
* The software supplied herewith by Microchip Technology Incorporated (the     *
* 'Company') is intended and supplied to you, the Company's customer, for use  *
* soley and exclusively on Microchip products.                                 *
*                                                                              *
* The software is owned by the Company and/or its supplier, and is protected   *
* under applicable copyright laws. All rights are reserved. Any use in         *
* violation of the foregoing restrictions may subject the user to criminal     *
* sanctions under applicable laws, as well as to civil liability for the       *
* breach of the terms and conditions of this license.                          *
*                                                                              *
* THIS SOFTWARE IS PROVIDED IN AN 'AS IS' CONDITION. NO WARRANTIES, WHETHER    *
* EXPRESS, IMPLIED OR STATUTORY, INCLUDING, BUT NOT LIMITED TO, IMPLIED        *
* WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE APPLY TO  *
* THIS SOFTWARE. THE COMPANY SHALL NOT, IN ANY CIRCUMSTANCES, BE LIABLE FOR    *
* SPECIAL, INCIDENTAL OR CONSEQUENTIAL DAMAGES, FOR ANY REASON WHATSOEVER.     *
********************************************************************************
*
* The following op-amps are covered by this model:
*      MCP606,MCP607,MCP608,MCP609
*
* Revision History:
*   REV A: 30-Jun-99, Created model
*   REV B: 18-Jul-02, Improved model
*   REV C: 12-Sep-06, Added over temperature, improved output stage, 
*                     fixed overdrive recovery time
*   REV D: 27-Jul-07, Updated output impedance for better model stability w/cap load,
*                     fixed CMRR freq shift
*
* Recommendations:
*      Use PSPICE (other simulators may require translation)
*      For a quick, effective design, use a combination of: data sheet
*            specs, bench testing, and simulations with this macromodel
*      For high impedance circuits, set GMIN=100F in the .OPTIONS statement
*
* Supported:
*      Typical performance for temperature range (-40 to 125) degrees Celsius
*      DC, AC, Transient, and Noise analyses.
*      Most specs, including: offsets, DC PSRR, DC CMRR, input impedance,
*            open loop gain, voltage ranges, supply current, ... , etc.
*      Temperature effects for Ibias, Iquiescent, Iout short circuit 
*            current, Vsat on both rails, Slew Rate vs. Temp and P.S.
*
* Not Supported:
*      Chip Select (MCP608)
*      Some Variation in specs vs. Power Supply Voltage
*      Monte Carlo (Vos, Ib),Process variation  
*      Distortion (detailed non-linear behavior)
*      Behavior outside normal operating region
*
* Input Stage
V10  3 10 900M
R10 10 11 2.18MEG
R11 10 12 2.18MEG
G10 10 11 10 11 45.8U
G11 10 12 10 12 45.8U
C11 11 12 3P
C12  1  0 6P
E12 71 14 POLY(6) 20 0 21 0 22 0 23 0 26 0 27 0
+ 90U 9.5 9.5 6 6 1 1
G12 1 0 62 0 1m
M12 11 14 15 15 NMI L=2.00U W=42.0U; *Added L & W values
M14 12 2 15 15 NMI L=2.00U W=42.0U; *Added L & W values
G14 2 0 62 0 1m
C13 1 2 0.5P
C14  2  0 6.00P
I15 15 4 5.00U
V16 16 4 -300M
GD16 16 1 TABLE {V(16,1)} ((-100,-1p)(0,0)(1m,1u)(2m,1m)) 
V13 3 13 1.1
GD13 2 13 TABLE {V(2,13)} ((-100,-1p)(0,0)(1m,1u)(2m,1m)) 
R71  1  0 20.0E12
R72  2  0 20.0E12
R73  1  2 20.0E12
I80  1  2 320E-15
*
* Noise, PSRR, and CMRR
I20 21 20 423U
D20 20  0 DN1
D21  0 21 DN1
I22 22 23 1N
R22 22 0  1k
R23  0 23 1k
G26  0 26 POLY(2) 3 0 4 0   0.00 -28.1U -3.5U
R26 26  0 1
G27  0 27 POLY(2) 1 0 2 0  -195U 11.2U 11.2U
R27 27  0 1
*
* Open Loop Gain, Slew Rate
G30  0 30 12 11 1
R30 30  0 1.00K
G31 0 31 3 4 0.00
I31 0 31 DC 91.3
R31 31  0 1 TC=2.60M,-7.26U
GD31 30 0 TABLE {V(30,31)} ((-100,-1n)(0,0)(1m,0.1)(2m,2))
G32 32 0 3 4 0.00
I32 32 0 DC 84
R32 32  0 1 TC=2.62M,-8.13U
GD32 0 30 TABLE {V(30,32)} ((-2m,2)(-1m,0.1)(0,0)(100,-1n))
G33  0 33 30 0 1m
R33  33 0 1K
G34  0 34 33 0 1.00
R34  34 0 1K
C34  34 0 950U
G37  0 37 34 0 1m
R37  37 0 1K
C37  37 0 1N
G371  0 371 37 0 1m
R371  371 0 1K
C371  371 0 100P
G38  0 38 371 0 1m 
R38  39 0 1K
L38  38 39 1.4M
E38  35 0 38 0 1
G35 33 0 TABLE {V(35,3)} ((-1,-1n)(0,0)(80,1n))(81,1))
G36 33 0 TABLE {V(35,4)} ((-81,-1)((-80,-1n)(0,0)(1,1n))
*
* Output Stage
R80 50 0 100MEG
G50 0 50 57 96 2
R58 57  96 0.50
R57 57  0 4.2k
C58  5  0 2.00P
G57  0 57 POLY(3) 3 0 4 0 35 0   0 0.145M 0.14M 0.3M
GD55 55 57 TABLE {V(55,57)} ((-2m,-1)(-1m,-1m)(0,0)(10,1n))
GD56 57 56 TABLE {V(57,56)} ((-2m,-1)(-1m,-1m)(0,0)(10,1n))
E55 55  0 POLY(2) 3 0 51 0 -1.6M 1 -32M
E56 56  0 POLY(2) 4 0 52 0 0.9M 1 -27M
R51 51 0 1k
R52 52 0 1k
GD51 50 51 TABLE {V(50,51)} ((-10,-1n)(0,0)(1m,1m)(2m,1))
GD52 50 52 TABLE {V(50,52)}  ((-2m,-1)(-1m,-1m)(0,0)(10,1n))
G53  3  0 POLY(1) 51 0  -5.00U 1M
G54  0  4 POLY(1) 52 0  -5.00U -1M
*
* Current Limit
G99 96 5 99 0 1
R98 0 98 1 TC=-4.46M,25.3U
G97 0 98 TABLE { V(96,5) } ((-11,-9.2M)(-1M,-9.1M)(0,0)(1M,9.1M)(11,9.2M))
E97 99 0 VALUE { V(98)*((V(3)-V(4))*293M + 266M)}
D98 4 5 DESD
D99 5 3 DESD
*
* Temperature / Voltage Sensitive IQuiscent
R61 0 61 1 TC=1.79M,-7.31U
G61 3 4 61 0 1
G60 0 61 TABLE {V(3, 4)} 
+ ((0,0)(900M,163N)(1.00,3.2U)(1.2,10.0U)
+ (1.6,11.1U)(2.2,16.3U)(5.5,18.6U))
*
* Temperature Sensitive offset voltage
I73 0 70 DC 1uA
R74 0 70 1 TC=-1.2,-75M
E75 1 71 70 0 1 
*
* Temp Sensistive IBias
I62 0 62 DC 1uA
R62 0 62 REXP  374.59883U
*
* Models
.MODEL NMI NMOS(KP=20.0U LEVEL=1 ); *Removed L & W values
.MODEL DESD  D   N=1 IS=1.00E-15
.MODEL DN1 D   IS=1P KF=.150F AF=1
.MODEL REXP RES TCE= 8.40918
.ENDS MCP606
