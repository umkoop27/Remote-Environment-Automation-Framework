.SUBCKT MCP616 1 2 3 4 5
*              | | | | |
*              | | | | Output
*              | | | Negative Supply
*              | | Positive Supply
*              | Inverting Input
*              Non-inverting Input
*
********************************************************************************
* Software License Agreement                                                   *
*                                                                              *
* The software supplied herewith by Microchip Technology Incorporated (the     *
* 'Company') is intended and supplied to you, the Company's customer, for use  *
* soley and exclusively on Microchip products.                                 *
*                                                                              *
* The software is owned by the Company and/or its supplier, and is protected   *
* under applicable copyright laws. All rights are reserved. Any use in         *
* violation of the foregoing restrictions may subject the user to criminal     *
* sanctions under applicable laws, as well as to civil liability for the       *
* breach of the terms and conditions of this license.                          *
*                                                                              *
* THIS SOFTWARE IS PROVIDED IN AN 'AS IS' CONDITION. NO WARRANTIES, WHETHER    *
* EXPRESS, IMPLIED OR STATUTORY, INCLUDING, BUT NOT LIMITED TO, IMPLIED        *
* WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE APPLY TO  *
* THIS SOFTWARE. THE COMPANY SHALL NOT, IN ANY CIRCUMSTANCES, BE LIABLE FOR    *
* SPECIAL, INCIDENTAL OR CONSEQUENTIAL DAMAGES, FOR ANY REASON WHATSOEVER.     *
********************************************************************************
*
* The following op-amps are covered by this model:
*      MCP616, MCP617, MCP618, MCP619
*
* Revision History:
*   REV A: 23-Feb-01, Created model
*   REV B: 19-Jul-02, Improved model 
*   REV C: 13-Sep-06, Added over temperature, improved output stage, 
*                     fixed overdrive recovery time
*   REV D: 27-Jul-07, Updated output impedance for better model stability w/cap load
*
* Recommendations:
*      Use PSPICE (other simulators may require translation)
*      For a quick, effective design, use a combination of: data sheet
*            specs, bench testing, and simulations with this macromodel
*      For high impedance circuits, set GMIN=100F in the .OPTIONS statement
*
* Supported:
*      Typical performance for temperature range (-40 to 125) degrees Celsius
*      DC, AC, Transient, and Noise analyses.
*      Most specs, including: offsets, DC PSRR, DC CMRR, input impedance,
*            open loop gain, voltage ranges, supply current, ... , etc.
*      Temperature effects for Ibias, Iquiescent, Iout short circuit 
*            current, Vsat on both rails, Slew Rate vs. Temp and P.S.
*
* Not Supported:
*      Chip Select (MCP618)
*      Some Variation in specs vs. Power Supply Voltage
*      Monte Carlo (Vos, Ib), Process variation
*      Distortion (detailed non-linear behavior)
*      Behavior outside normal operating region
*
* Input Stage
V10  3 10 0.68
R10 10 11 1.54MEG
R11 10 12 1.54MEG
G10 10 11 10 11 64.8U
G11 10 12 10 12 64.8U
C11 11 12 12P
C12  1  0 3.70P
E12 71 14 POLY(6) 20 0 21 0 22 0 23 0 26 0 27 0
+ 120U 6.85 6.85 4.2 4.2 1 1
G12 1 0 62 0 -1m
G13 1 2 63 0 1m
M12 11 14 15 15 NMI L=2.00U W=42.0U; *Added L & W values
M14 12 2 15 15 NMI L=2.00U W=42.0U; *Added L & W values
G14 2 0 62 0 -1m
C14  2  0 3.70P
I15 15 4 10.0U
V16 16 4 -10m
GD16 16 1 TABLE {V(16,1)} ((-100,-1p)(0,0)(1m,1u)(2m,1m)) 
V13 3 13 880M
GD13 2 13 TABLE {V(2,13)} ((-100,-1p)(0,0)(1m,1u)(2m,1m)) 
R71  1  0 600MEG
R72  2  0 600MEG
R73  1  2 3.00MEG
I80  1  2 75.0P
*
* Noise, PSRR, and CMRR
I20 21 20 423U
D20 20  0 DN1
D21  0 21 DN1
I22 22 23 1N
R22 22 0  1k
R23  0 23 1k
G26  0 26 POLY(2) 3 0 4 0   0.00 -2.2U -6.2U
R26 26  0 1
G27  0 27 POLY(2) 1 0 2 0  -61.7U 3U 3U
R27 27  0 1
*
* Open Loop Gain, Slew Rate
G30  0 30 12 11 1
R30 30  0 1K
G31 0 31 3 4 0.00
I31 0 31 DC 64.0
R31 31  0 1.06 TC=2.2M,-1U
GD31 30 0 TABLE {V(30,31)} ((-100,-1n)(0,0)(1m,0.1)(2m,2))
G32 32 0 3 4 0.00
I32 32 0 DC 53.8
R32 32  0 1.06 TC=2.3M,-1U
GD32 0 30 TABLE {V(30,32)} ((-2m,2)(-1m,0.1)(0,0)(100,-1n))
G33  0 33 30 0 1m
R33  33 0 1K
G34  0 34 33 0 1.77
R34  34 0 1K
C34  34 0 1.49M
G37  0 37 34 0 1m
R37  37 0 1K
C37  37 0 1.8N
G371  0 371 37 0 1m
R371  371 0 1K
C371  371 0 62P
G38  0 38 371 0 1m
R38  39 0 1K
L38  38 39 1.8M
E38  35 0 38 0 1
G35 33 0 TABLE {V(35,3)} ((-1,-1n)(0,0)(120,1n))(121,1))
G36 33 0 TABLE {V(35,4)} ((-121,-1)((-120,-1n)(0,0)(1,1n))
*
* Output Stage
R80 50 0 100MEG
G50 0 50 57 96 2
R58 57  96 0.50
R57 57  0 5000
C58  5  0 2.00P
G57  0 57 POLY(3) 3 0 4 0 35 0   0 75U 75U 200U
GD55 55 57 TABLE {V(55,57)} ((-2m,-1)(-1m,-1m)(0,0)(10,1n))
GD56 57 56 TABLE {V(57,56)} ((-2m,-1)(-1m,-1m)(0,0)(10,1n))
E55 55  0 POLY(2) 3 0 51 0 -0.7M 1 -61.1M
E56 56  0 POLY(2) 4 0 52 0 1M 1 -51.3M
R51 51 0 1k
R52 52 0 1k
GD51 50 51 TABLE {V(50,51)} ((-10,-1n)(0,0)(1m,1m)(2m,1))
GD52 50 52 TABLE {V(50,52)}  ((-2m,-1)(-1m,-1m)(0,0)(10,1n))
G53  3  0 POLY(1) 51 0  -9.65U 1M
G54  0  4 POLY(1) 52 0  -9.65U -1M
*
* Current Limit
G99 96 5 99 0 1
R98 0 98 1 TC=-5.41M,11.3U
G97 0 98 TABLE { V(96,5) } ((-11.0,-8.7M)(-1.00M,-8.61M)(0,0)(1.00M,8.61M)(11.0,8.7M))
E97 99 0 VALUE { V(98)*((V(3)-V(4))*298M + 314M)}
D98 4 5 DESD
D99 5 3 DESD
*
* Temperature / Voltage Sensitive IQuiscent
R61 0 61 1 TC=3.0M,-3U
G61 3 4 61 0 1
G60 0 61 TABLE {V(3, 4)} 
+ ((0,0)(800M,10N)(1.3,13.2U)(1.5,14.3U)
+ (1.6,13.9U)(2.1,17.4U)(5.5,19.4U))
*
* Temperature Sensitive offset voltage
I73 0 70 DC 1uA
R74 0 70 1 TC=2.5
E75 1 71 70 0 1 
*
* Temp Sensistive IBias
I62 0 62 DC 1uA
R62 0 62 16.6 TC=-4.5M,20U
I63 0 63 DC 1uA
R63 0 63 180m TC=-16.4M,25U
*
* Models
.MODEL NMI NMOS(KP=20.0U LEVEL=1 ); *Removed L * W values
.MODEL DESD  D   N=1 IS=1.00E-15
.MODEL DN1 D   IS=1P KF=146E-18 AF=1
.ENDS MCP616
