.SUBCKT MCP6V01 1 2 3 4 5
*               | | | | |
*               | | | | Output
*               | | | Negative Supply
*               | | Positive Supply
*               | Inverting Input
*               Non-inverting Input
*
********************************************************************************
* Software License Agreement                                                   *
*                                                                              *
* The software supplied herewith by Microchip Technology Incorporated (the     *
* 'Company') is intended and supplied to you, the Company's customer, for use  *
* soley and exclusively on Microchip products.                                 *
*                                                                              *
* The software is owned by the Company and/or its supplier, and is protected   *
* under applicable copyright laws. All rights are reserved. Any use in         *
* violation of the foregoing restrictions may subject the user to criminal     *
* sanctions under applicable laws, as well as to civil liability for the       *
* breach of the terms and conditions of this license.                          *
*                                                                              *
* THIS SOFTWARE IS PROVIDED IN AN 'AS IS' CONDITION. NO WARRANTIES, WHETHER    *
* EXPRESS, IMPLIED OR STATUTORY, INCLUDING, BUT NOT LIMITED TO, IMPLIED        *
* WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE APPLY TO  *
* THIS SOFTWARE. THE COMPANY SHALL NOT, IN ANY CIRCUMSTANCES, BE LIABLE FOR    *
* SPECIAL, INCIDENTAL OR CONSEQUENTIAL DAMAGES, FOR ANY REASON WHATSOEVER.     *
********************************************************************************
*
* The following op-amps are covered by this model:
*      MCP6V01, MCP6V02, MCP6V03
*
* Revision History:
*      REV A: 9/15/2008, Created model
*      REV B: 8/15/2009, fixed the output swing issue for voltage follower application
*
* Recommendations:
*      Use PSPICE (or SPICE 2G6; other simulators may require translation)
*      For a quick, effective design, use a combination of: data sheet
*            specs, bench testing, and simulations with this macromodel
*      For high impedance circuits, set GMIN=100F in the .OPTIONS statement
*
* Supported:
*      Typical performance for temperature range (-40 to 125) degrees Celsius
*      DC, AC, Transient, and Noise analyses.
*      Most specs, including: offsets, DC PSRR, DC CMRR, input impedance,
*            open loop gain, voltage ranges, supply current, ... , etc.
*      Temperature effects for Ibias, Iquiescent, Iout short circuit 
*            current, Vsat on both rails, Slew Rate vs. Temp and P.S.
*
* Not Supported:
*      Some Variation in specs vs. Power Supply Voltage
*      Monte Carlo (Vos, Ib), Process variation
*      Distortion (detailed non-linear behavior)
*      Some Temperature analysis
*      Behavior outside normal operating region
*
* Input Stage
V10  3 10 -400M
R10 10 11 690K
R11 10 12 690K
G10 10 11 10 11 144U
G11 10 12 10 12 144U
C11 11 12 0.8P
C12  1  0 6P
E12 71 14 POLY(4) 200 0 220 0 26 0 27 0 -1u 5 20 1 1
G12 1 0 62 0 1m
G13 1 2 63 0 1u
M12 11 14 15 15 NMI L=2.00U W=42.0U; *Added L & W values
M14 12 2 15 15 NMI L=2.00U W=42.0U; *Added L & W values
G14 2 0 62 0 1m
C13  1  2 3P
C14  2  0 6P
I15 15 4 50U
V16 16 4 -200m
GD16 16 1 TABLE {V(16,1)} ((-100,-1p)(0,0)(1m,1u)(2m,1m)) 
V13 3 13 -200m
GD13 2 13 TABLE {V(2,13)} ((-100,-1p)(0,0)(1m,1u)(2m,1m))
R71  1  0 11T
R72  2  0 11T
R73  1  2 11T
*
* Noise, PSRR, and CMRR
I20 21 20 423U
D20 20  0 DN1
D21  0 21 DN1
G20 200 0 POLY(2) 21 0 20 0 0 1m 1m
R20 200 0 1k
I22 22 23 1N
R22 22 0  1k
R23  0 23 1k
G22 220 0 POLY(2) 22 0 23 0 0 1m 1m
R220 220 0 1k
R221 220 221 400
C221 221 0 20N
G26  0 26 POLY(2) 3 0 4 0   0.00 -40N -40N
R26 26  0 1
G27  0 27 POLY(2) 1 0 2 0  -1.73U 20N 20N
R27 27  0 1
*These statements will put in correct CMRR curve over 1MHz, but slows simulation slightly and R271 increases noise above 50kHz
*R27 27  271 1
*L27 271  0 500m
*R271 271 0 0.7MEG
*C27 271  0 0.5p
*
* Open Loop Gain, Slew Rate
G30  0 30 12 11 1
R30 30  0 1.00K
G31 0 31 3 4 4.5
I31 0 31 DC 19
R31 31  0 1 TC=1.43M, -2U
GD31 30 0 TABLE {V(30,31)} ((-100,-1n)(0,0)(1m,0.1)(2m,2))
G32 32 0 3 4 -0.5
I32 32 0 DC 40
R32 32  0 1 TC=1.07M,-2.36U
GD32 0 30 TABLE {V(30,32)} ((-2m,2)(-1m,0.1)(0,0)(100,-1n))
G33  0 33 30 0 1m
R33  33 0 1K
G34  0 34 33 0 50
R34  34 0 1K
C34  34 0 2.5M
G37  0 37 34 0 1m
R37  37 0 1K
C37  37 371 120P
RC37 371 0 100
G38  0 38 37 0 1m
R38  39 0 1K
L38  38 39 220U
E38  35 0 38 0 1
G35 33 0 TABLE {V(35,3)} ((-1,-1n)(0,0)(25.0,1n))(26,1))
G36 33 0 TABLE {V(35,4)} ((-18,-1)((-17,-1n)(0,0)(1,1n))
*
* Output Stage
R80 50 0 100MEG
G50 0 50 57 96 1
R58 57  96 0.50
R57 57  0 1k
C58  5  0 2.00P
G57  0 57 POLY(3) 3 0 4 0 35 0   0 1.5M 1.3M 833U
GD55 55 57 TABLE {V(55,57)} ((-2m,-1)(-1m,-1m)(0,0)(10,1n))
GD56 57 56 TABLE {V(57,56)} ((-2m,-1)(-1m,-1m)(0,0)(10,1n))
E55 55  0 POLY(2) 3 0 51 0 -5M  1.002 -145M   0   25M    0
E56 56  0 POLY(2) 4 0 52 0 7M 1  -34M 0  10M  20M
R51 51 0 1k
R52 52 0 1k
GD51 50 51 TABLE {V(50,51)} ((-10,-1n)(0,0)(1m,1m)(2m,1))
GD52 50 52 TABLE {V(50,52)}  ((-2m,-1)(-1m,-1m)(0,0)(10,1n))
G53  3  0 POLY(1) 51 0  -50.0U 1M
G54  0  4 POLY(1) 52 0  -50.0U -1M
*
* Current Limit
G99 96 5 99 0 1
R98 0 98 1 TC=-4.86M,26.4U
G97 0 98 TABLE { V(96,5) } ((-11,-9M)(-1M,-8.91M)(0,0)(1M,9.91M)(11,10M))
E97 99 0 VALUE { V(98)*((V(3)-V(4))*355M + 288M)}
D98 4 5 DESD
D99 5 3 DESD
*
* Temperature / Voltage Sensitive IQuiscent
R61 0 61 1 TC=1.86M,-3.01U
G61 3 4 61 0 1
G60 0 61 TABLE {V(3, 4)} 
+ ((0,0)(900M,3.25U)(1.4,260U)(1.5,280U)
+ (3.5,300U)(5.5,325U)(6.5,355U))
*
* Temperature Sensitive offset voltage
I73 0 70 DC 1uA
R74 0 70 1 TC=50.0M
E75 1 71 70 0 1 
*
* Temp Sensistive IBias
I62 0 62 DC 1uA
R62 0 62 REXP  2.03M
*
* Temp Sensistive Offset IBias
I63 0 63 DC 1uA
R63 0 63 15 TC=-2M,180U
*
* Models
.MODEL NMI NMOS(KP=20.0U LEVEL=1 ); *Removed L & W values
.MODEL DESD  D   N=2 IS=1.00E-15
.MODEL DN1 D   IS=1P KF=146E-18 AF=1
.MODEL REXP  RES TCE= 5.86758
.ENDS MCP6V01
